* /home/sumanto/Desktop/verilog/eSim/One_Hot_Counter/One_Hot_Counter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun Nov 21 19:26:26 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_U2-Pad1_ GND pulse		
v2  Net-_U2-Pad2_ GND pulse		
v3  Net-_U2-Pad3_ GND pulse		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ adc_bridge_3		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ ? ? ? ? ? ? ? ? one_hot_cnt		

.end
