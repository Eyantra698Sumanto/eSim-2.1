* /home/sumanto/Desktop/verilog/eSim/i2c/i2c.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun Nov 21 23:55:39 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U4  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ Net-_U2-Pad10_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ Net-_U3-Pad13_ Net-_U3-Pad14_ ? ? ? ? ? ? ? ? ? ? ? ? ? ? i2c_master_top		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ counter3bit		
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ Net-_U2-Pad9_ Net-_U2-Pad10_ counter8bit		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U3-Pad3_ Net-_U3-Pad4_ Net-_U3-Pad5_ Net-_U3-Pad6_ Net-_U3-Pad7_ Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U3-Pad10_ Net-_U3-Pad11_ Net-_U3-Pad12_ Net-_U3-Pad13_ Net-_U3-Pad14_ adc_bridge_7		
v4  Net-_U3-Pad4_ GND pulse		
v5  Net-_U3-Pad5_ GND pulse		
v6  Net-_U3-Pad6_ GND pulse		
v7  Net-_U3-Pad7_ GND pulse		
v3  Net-_U3-Pad3_ GND pulse		
v2  Net-_U3-Pad2_ GND pulse		
v1  Net-_U3-Pad1_ GND pulse		

.end
