/* verilator lint_off UNUSED */
module hello;
////fvcgg
///hello
//good good
//oh!
//jggjgj
//f
//Sumanto
initial
    begin
    $display("Hello world");
    $finish;
    end
endmodule
