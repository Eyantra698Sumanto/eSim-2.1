* /home/sumanto/Desktop/verilog/eSim/interruptcontroller/interruptcontroller.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue Nov 30 10:16:57 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U10-Pad6_ Net-_U10-Pad7_ Net-_U10-Pad8_ Net-_U10-Pad9_ Net-_U10-Pad10_ counter8bit		
v1  clk GND pulse		
v2  rst GND pulse		
v3  intr_in GND pulse		
U5  clk rst intr_in Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad19_ adc_bridge_3		
U1  clk plot_v1		
U2  rst plot_v1		
U4  intr_in plot_v1		
U7  Net-_U10-Pad20_ Net-_U10-Pad21_ intr_out busoe dac_bridge_2		
U8  intr_out plot_v1		
U9  busoe plot_v1		
U10  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad3_ Net-_U10-Pad4_ Net-_U10-Pad5_ Net-_U10-Pad6_ Net-_U10-Pad7_ Net-_U10-Pad8_ Net-_U10-Pad9_ Net-_U10-Pad10_ Net-_U10-Pad11_ Net-_U10-Pad12_ Net-_U10-Pad13_ Net-_U10-Pad14_ Net-_U10-Pad15_ Net-_U10-Pad16_ Net-_U10-Pad17_ Net-_U10-Pad18_ Net-_U10-Pad19_ Net-_U10-Pad20_ Net-_U10-Pad21_ intr_cntrl		
U6  Net-_U10-Pad1_ Net-_U10-Pad2_ Net-_U10-Pad11_ Net-_U10-Pad12_ Net-_U10-Pad13_ Net-_U10-Pad14_ Net-_U10-Pad15_ Net-_U10-Pad16_ Net-_U10-Pad17_ Net-_U10-Pad18_ counter8bit		

.end
