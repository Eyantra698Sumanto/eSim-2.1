* /home/sumanto/Desktop/verilog/eSim/calculator/calculator.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Nov 29 00:59:18 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U1-Pad18_ ? ? ? ? ? ? ? ? ? ? ? calculator		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ ? ? Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U1-Pad11_ Net-_U1-Pad12_ Net-_U1-Pad13_ Net-_U1-Pad14_ Net-_U1-Pad15_ Net-_U1-Pad16_ Net-_U1-Pad17_ Net-_U1-Pad18_ counter16bit		
U3  Net-_U3-Pad1_ Net-_U3-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
v1  Net-_U3-Pad1_ GND pulse		
v2  Net-_U3-Pad2_ GND pulse		

.end
