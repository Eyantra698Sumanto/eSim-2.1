* /home/sumanto/Desktop/verilog/eSim/microcomputer/microcomputer.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Nov 22 01:31:32 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? cpu		
v1  Net-_U2-Pad1_ GND pulse		
U2  Net-_U2-Pad1_ Net-_U1-Pad1_ adc_bridge_1		

.end
