* /home/sumanto/Desktop/verilog/eSim/parallel_crc/parallel_crc.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun Nov 21 15:25:50 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U3  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? ? parallel_crc		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ counter8bit		
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_4		
v1  Net-_U2-Pad1_ GND pulse		
v2  Net-_U2-Pad2_ GND pulse		
v3  Net-_U2-Pad3_ GND pulse		
v4  Net-_U2-Pad4_ GND pulse		

.end
