* /home/sumanto/Desktop/verilog/eSim/basicgates/basicgates.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Nov  8 16:16:55 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ jbasicgates		
U4  A B Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
U5  Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U2-Pad7_ Net-_U2-Pad8_ OROUT ANDOUT XOR NOR NAND XNOR dac_bridge_6		
v1  A GND pulse		
v2  B GND pulse		
U1  A plot_v1		
U3  B plot_v1		
U6  OROUT plot_v1		
U7  ANDOUT plot_v1		
U8  XOR plot_v1		
U9  NOR plot_v1		
U10  NAND plot_v1		
U11  XNOR plot_v1		

.end
