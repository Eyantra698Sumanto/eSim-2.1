
/* verilator lint_off UNUSED */
/* verilator lint_off EOFNEWLINE */
/* verilator lint_off DECLFILENAME */
/* verilator lint_off BLKSEQ */
/* verilator lint_off WIDTH */
/* verilator lint_off LATCH */
/* verilator lint_off SELRANGE */
/* verilator lint_off PINCONNECTEMPTY */
/* verilator lint_off DEFPARAM */
/* verilator lint_off IMPLICIT */
/* verilator lint_off TIMESCALEMOD */
/* verilator lint_off COMBDLY */
/* verilator lint_off SYNCASYNCNET */
/* verilator lint_off UNOPTFLAT */
/* verilator lint_off UNSIGNED */
/* verilator lint_off CASEINCOMPLETE */
/* verilator lint_off UNDRIVEN */
    `line 2 "trafficmaker.tlv" 0 //_\TLV_version 1d: tl-x.org, generated by SandPiper(TM) 1.11-2021/01/28-beta
`include "sp_default.vh" //_\SV
                 
//_\SV
   module trafficmaker(input wire clk, input wire reset, input wire [31:0] cyc_cnt, output wire passed, output wire failed);    /* verilator lint_save */ /* verilator lint_off UNOPTFLAT */  bit [256:0] RW_rand_raw; bit [256+63:0] RW_rand_vect; pseudo_rand #(.WIDTH(257)) pseudo_rand (clk, reset, RW_rand_raw[256:0]); assign RW_rand_vect[256+63:0] = {RW_rand_raw[62:0], RW_rand_raw};  /* verilator lint_restore */  /* verilator lint_off WIDTH */ /* verilator lint_off UNOPTFLAT */  
   //BY SUMANTO KAR
   wire [15:0] led;
   reg [3:0] digit;
   reg [6:0] segment;
   wire  dp = 1;
 
   reg [2:0] state;
   reg [2:0] count;
 
   parameter [2:0] NORTH    =   3'b000;
   parameter [2:0] NORTH_Y  =   3'b001;
   parameter [2:0] SOUTH    =   3'b010;
   parameter [2:0] SOUTH_Y  =   3'b011;
   parameter [2:0] EAST     =   3'b100;
   parameter [2:0] EAST_Y   =   3'b101;
   parameter [2:0] WEST     =   3'b110;
   parameter [2:0] WEST_Y   =   3'b111;

   always @(posedge clk, posedge reset)
     begin
        if (reset)
            begin
               assign state=NORTH;
               assign count=3'b000;
               
                /* TODO: Set initial state to NORTH and count signal to zero */
                // 
                // 
               
            end
        else
            begin
                case (state)
                NORTH :
                    begin
                       
                       // Enable first seven segment and set to Green 
                       digit <= 4'b0111;
                       segment <= 7'b1110111;
                       
                        /* TODO: 1. Keep the green NORTH signal active for 8 seconds 
                                2. Set state of signal to yellow NORTH after that 
                          HINT: Use if-else block
                        */
                       if(count==7) begin
                             assign state=NORTH_Y;
                              assign count=0;    
                          end
                       else assign count=count+1;
                                                  
                             
                       
                    end

                NORTH_Y :
                    begin
                       
                        // Enable first seven segment and set to Yellow
                        digit <= 4'b0111;
                        segment <= 7'b1111110;
                       
                        /* TODO: 1. Keep the yellow NORTH signal active for 4 seconds 
                                2. Set state of signal to green SOUTH after that 
                        */
                      if(count==3) begin
                             assign state=SOUTH;
                              assign count=0;    
                          end
                       else assign count=count+1;
                            end
               SOUTH :
                    begin
                       
                        // TODO: Enable second seven segment and set to Green 
                       digit <= 4'b1011;
                       segment <= 7'b1110111;
                        /* TODO: 1. Keep the green SOUTH signal active for 8 seconds 
                                 2. Set state of signal to yellow SOUTH after that 
                        */
                       if(count==7) begin
                             assign state=SOUTH_Y;
                              assign count=0;    
                          end
                       else assign count=count+1;
                    end

                SOUTH_Y :
                    begin
                    
                        // TODO: Enable second seven segment and set to Yellow 
                            digit <= 4'b1011;
                        segment <= 7'b1111110;
                        /* TODO: 1. Keep the yellow SOUTH signal active for 4 seconds 
                                    2. Set state of signal to green EAST after that 
                        */
                    if(count==3) begin
                             assign state=EAST;
                              assign count=0;    
                          end
                       else assign count=count+1;
                   end
                EAST :
                    begin
                       
                    
                        // TODO: Enable third seven segment and set to Green 
                            digit <= 4'b1101;
                        segment <= 7'b1110111;
                        /* TODO: 1. Keep the green EAST signal active for 8 seconds 
                                2. Set state of signal to yellow EAST after that 
                        */
                       if(count==7) begin
                             assign state=EAST_Y;
                              assign count=0;    
                          end
                       else assign count=count+1;
                    
                    end
                EAST_Y :
                    begin
                    
                    // TODO: Enable third seven segment and set to Yellow 
                    digit <= 4'b1101;
                    segment <= 7'b1111110;
                    /* TODO: 1. Keep the yellow EAST signal active for 4 seconds 
                                2. Set state of signal to green WEST after that 
                    */
                          if(count==3) begin
                             assign state=WEST;
                              assign count=0;    
                          end
                       else assign count=count+1;
                    end
                WEST :
                    begin

                    // TODO: Enable fourth seven segment and set to Green 
                            digit <= 4'b1110;
                       segment <= 7'b1110111;
                    /* TODO: 1. Keep the green WEST signal active for 8 seconds 
                            2. Set state of signal to yellow WEST after that 
                    */
                            if(count==7) begin
                             assign state=WEST_Y;
                              assign count=0;    
                          end
                       else assign count=count+1;
                    end
                WEST_Y :
                    begin

                    // TODO: Enable fourth seven segment and set to Yellow 
                            digit <= 4'b1110;
                     segment <= 7'b1111110;
                    /* TODO: 1. Keep the yellow EAST signal active for 4 seconds 
                            2. Move back to NORTH signal again
                    */
                            if(count==3) begin
                             assign state=NORTH;
                              assign count=0;    
                          end
                       else assign count=count+1;
                    end
                 
            endcase 
        end 
    end 
    assign led = count;

`include "trafficmaker_gen.sv" //_\TLV
   // M4_BOARD numbering
   // 1 - Zedboard
   // 2 - Artix-7
   // 3 - Basys3
   // 4 - Icebreaker
   // 5 - Nexys
   
   `line 33 "fpgaincludes.tlv" 1   // Instantiated from trafficmaker.tlv, 184 as: m4+fpga_init()
      //m4+osfpga_logo()
      //_|fpga_init_macro
         //_@0
            
            
            
               
                     
                     
                           
                           
                              
                              
                           
                           
                            
                            
                            
                            
                            
                            
                           
                        
                   
            
            
            
               
                     
                     
                           
                           
                              
                              
                           
                           
                            
                            
                            
                            
                            
                            
                           
                        
                     
                        
                        
                        
                        
                        
                        
                     
                   
                   
                   
            
               
                  
                     
                        
                              
                              
                              
                              
                              
                           
                           
                           
                              
                              
                              
                              
                              
                              
                              
                           
                        
                     
            
            
            
               
                     
                     
                           
                           
                              
                              
                           
                           
                            
                            
                            
                            
                            
                            
                           
                        
                     
                              
                              
                              
                              
                              
                              
                           
                   
                   
            
               
                  
                     
                        
                              
                              
                              
                              
                              
                           
                           
                           
                              
                              
                              
                              
                              
                              
                              
                           
                        
                     
            
            
            
               
                     
                     
                     
                           
                           
                              
                              
                           
                           
                            
                            
                            
                            
                            
                            
                           
                        
                   
            
            
            
               
                     
                     
                           
                           
                              
                              
                           
                           
                            
                            
                            
                           
                        
                   
                        
                        
                        
                        
                        
                        
                     
                   
                   
                
            
               
                  
                     
                        
                              
                              
                              
                              
                              
                              
                           
                           
                           
                              
                              
                              
                              
                              
                              
                              
                           
                        
                     
            
            
            
            
            
            
            
   //_\end_source
   `line 185 "trafficmaker.tlv" 2
   `line 246 "fpgaincludes.tlv" 1   // Instantiated from trafficmaker.tlv, 185 as: m4+fpga_led(*led)
      //_|led_pipe_macro
         //_@0
            
            
            
            
               
                  
                     
                           
                           
                           
                           
                           
                           
                        
                     
                  
                  
                        
                        
                     
            
            
            
               
                  
                     
                           
                           
                           
                           
                           
                           
                        
                     
                  
                  
                        
                        
                     
            
            
            
               
                  
                     
                           
                           
                           
                           
                           
                           
                        
                     
                  
                  
                        
                        
                     
            
            
   
            
            
            
            
               
                  
                     
                           
                           
                           
                           
                           
                           
                        
                     
                  
                  
                        
                        
                  
            
            
            
            
            
            
            
   //_\end_source
   `line 186 "trafficmaker.tlv" 2
   `line 357 "fpgaincludes.tlv" 1   // Instantiated from trafficmaker.tlv, 186 as: m4+fpga_sseg(*digit, *segment, *dp)
      //_|sseg_pipe_macro
         //_@0
            
            
            
            
            
            
            
            
               
                  
                     
                        
                              
                              
                              
                              
                              
                           
                           
                           
                              
                              
                              
                              
                              
                              
                              
                           
                        
                     
                     
                        
                        
                        
                        
                        
                           
                        
                        
                           
                           
                        
                     
            
            
            
               
                  
                     
                        
                              
                              
                              
                              
                              
                           
                           
                           
                              
                              
                              
                              
                              
                              
                              
                           
                        
                     
                     
                        
                        
                        
                        
                        
                           
                        
                        
                           
                           
                        
                     
            
            
            
               
                  
                  
                        
                        
                           
                           
                        
                        
                         
                         
                         
                         
                         
                        
                     
                   
                        
                        
                           
                           
                        
                        
                         
                         
                         
                         
                         
                        
                     
                   
                     
                     
                     
                     
                     
                     
                  
                  
                     
                     
                     
                     
                     
                     
                  
                
                
            
               
                  
                     
                        
                              
                              
                              
                              
                              
                           
                           
                           
                              
                              
                              
                              
                              
                              
                              
                           
                        
                     
                     
                        
                        
                        
                        
                        
                        
                           
                        
                        
                           
                           
                        
                     
            
            
            
               
                  
                     
                        
                              
                              
                              
                              
                              
                              
                           
                           
                           
                              
                              
                              
                              
                              
                              
                              
                           
                        
                     
                     
                        
                        
                        
                        
                        
                           
                        
                        
                           
                           
                        
                     
            
            
            
            
            
            
   //_\end_source
   `line 187 "trafficmaker.tlv" 2
   assign passed = led > 6; endgenerate
//_\SV
   endmodule

