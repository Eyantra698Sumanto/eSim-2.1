* /home/sumanto/Desktop/verilog/eSim/xorxnor/xorxnor.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Thu Nov 11 00:28:49 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ ixorxnor		
U4  A B Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U5  Net-_U1-Pad3_ Net-_U1-Pad4_ XOR XNOR dac_bridge_2		
v1  A GND pulse		
v2  B GND pulse		
U2  A plot_v1		
U3  B plot_v1		
U6  XOR plot_v1		
U7  XNOR plot_v1		

.end
