
/* verilator lint_off UNUSED */
/* verilator lint_off EOFNEWLINE */
/* verilator lint_off DECLFILENAME */
/* verilator lint_off BLKSEQ */
/* verilator lint_off WIDTH */
/* verilator lint_off LATCH */
/* verilator lint_off SELRANGE */
/* verilator lint_off PINCONNECTEMPTY */
/* verilator lint_off DEFPARAM */
/* verilator lint_off IMPLICIT */
/* verilator lint_off TIMESCALEMOD */
/* verilator lint_off COMBDLY */
/* verilator lint_off SYNCASYNCNET */
/* verilator lint_off UNOPTFLAT */
    module aes_sbox(ip,op);
input	[7:0]	ip;
output	[7:0]	op;
reg	[7:0]	op;

always @(ip)
	case(ip)		
	   8'h00: op=8'h63;
	   8'h01: op=8'h7c;
	   8'h02: op=8'h77;
	   8'h03: op=8'h7b;
	   8'h04: op=8'hf2;
	   8'h05: op=8'h6b;
	   8'h06: op=8'h6f;
	   8'h07: op=8'hc5;
	   8'h08: op=8'h30;
	   8'h09: op=8'h01;
	   8'h0a: op=8'h67;
	   8'h0b: op=8'h2b;
	   8'h0c: op=8'hfe;
	   8'h0d: op=8'hd7;
	   8'h0e: op=8'hab;
	   8'h0f: op=8'h76;
	   8'h10: op=8'hca;
	   8'h11: op=8'h82;
	   8'h12: op=8'hc9;
	   8'h13: op=8'h7d;
	   8'h14: op=8'hfa;
	   8'h15: op=8'h59;
	   8'h16: op=8'h47;
	   8'h17: op=8'hf0;
	   8'h18: op=8'had;
	   8'h19: op=8'hd4;
	   8'h1a: op=8'ha2;
	   8'h1b: op=8'haf;
	   8'h1c: op=8'h9c;
	   8'h1d: op=8'ha4;
	   8'h1e: op=8'h72;
	   8'h1f: op=8'hc0;
	   8'h20: op=8'hb7;
	   8'h21: op=8'hfd;
	   8'h22: op=8'h93;
	   8'h23: op=8'h26;
	   8'h24: op=8'h36;
	   8'h25: op=8'h3f;
	   8'h26: op=8'hf7;
	   8'h27: op=8'hcc;
	   8'h28: op=8'h34;
	   8'h29: op=8'ha5;
	   8'h2a: op=8'he5;
	   8'h2b: op=8'hf1;
	   8'h2c: op=8'h71;
	   8'h2d: op=8'hd8;
	   8'h2e: op=8'h31;
	   8'h2f: op=8'h15;
	   8'h30: op=8'h04;
	   8'h31: op=8'hc7;
	   8'h32: op=8'h23;
	   8'h33: op=8'hc3;
	   8'h34: op=8'h18;
	   8'h35: op=8'h96;
	   8'h36: op=8'h05;
	   8'h37: op=8'h9a;
	   8'h38: op=8'h07;
	   8'h39: op=8'h12;
	   8'h3a: op=8'h80;
	   8'h3b: op=8'he2;
	   8'h3c: op=8'heb;
	   8'h3d: op=8'h27;
	   8'h3e: op=8'hb2;
	   8'h3f: op=8'h75;
	   8'h40: op=8'h09;
	   8'h41: op=8'h83;
	   8'h42: op=8'h2c;
	   8'h43: op=8'h1a;
	   8'h44: op=8'h1b;
	   8'h45: op=8'h6e;
	   8'h46: op=8'h5a;
	   8'h47: op=8'ha0;
	   8'h48: op=8'h52;
	   8'h49: op=8'h3b;
	   8'h4a: op=8'hd6;
	   8'h4b: op=8'hb3;
	   8'h4c: op=8'h29;
	   8'h4d: op=8'he3;
	   8'h4e: op=8'h2f;
	   8'h4f: op=8'h84;
	   8'h50: op=8'h53;
	   8'h51: op=8'hd1;
	   8'h52: op=8'h00;
	   8'h53: op=8'hed;
	   8'h54: op=8'h20;
	   8'h55: op=8'hfc;
	   8'h56: op=8'hb1;
	   8'h57: op=8'h5b;
	   8'h58: op=8'h6a;
	   8'h59: op=8'hcb;
	   8'h5a: op=8'hbe;
	   8'h5b: op=8'h39;
	   8'h5c: op=8'h4a;
	   8'h5d: op=8'h4c;
	   8'h5e: op=8'h58;
	   8'h5f: op=8'hcf;
	   8'h60: op=8'hd0;
	   8'h61: op=8'hef;
	   8'h62: op=8'haa;
	   8'h63: op=8'hfb;
	   8'h64: op=8'h43;
	   8'h65: op=8'h4d;
	   8'h66: op=8'h33;
	   8'h67: op=8'h85;
	   8'h68: op=8'h45;
	   8'h69: op=8'hf9;
	   8'h6a: op=8'h02;
	   8'h6b: op=8'h7f;
	   8'h6c: op=8'h50;
	   8'h6d: op=8'h3c;
	   8'h6e: op=8'h9f;
	   8'h6f: op=8'ha8;
	   8'h70: op=8'h51;
	   8'h71: op=8'ha3;
	   8'h72: op=8'h40;
	   8'h73: op=8'h8f;
	   8'h74: op=8'h92;
	   8'h75: op=8'h9d;
	   8'h76: op=8'h38;
	   8'h77: op=8'hf5;
	   8'h78: op=8'hbc;
	   8'h79: op=8'hb6;
	   8'h7a: op=8'hda;
	   8'h7b: op=8'h21;
	   8'h7c: op=8'h10;
	   8'h7d: op=8'hff;
	   8'h7e: op=8'hf3;
	   8'h7f: op=8'hd2;
	   8'h80: op=8'hcd;
	   8'h81: op=8'h0c;
	   8'h82: op=8'h13;
	   8'h83: op=8'hec;
	   8'h84: op=8'h5f;
	   8'h85: op=8'h97;
	   8'h86: op=8'h44;
	   8'h87: op=8'h17;
	   8'h88: op=8'hc4;
	   8'h89: op=8'ha7;
	   8'h8a: op=8'h7e;
	   8'h8b: op=8'h3d;
	   8'h8c: op=8'h64;
	   8'h8d: op=8'h5d;
	   8'h8e: op=8'h19;
	   8'h8f: op=8'h73;
	   8'h90: op=8'h60;
	   8'h91: op=8'h81;
	   8'h92: op=8'h4f;
	   8'h93: op=8'hdc;
	   8'h94: op=8'h22;
	   8'h95: op=8'h2a;
	   8'h96: op=8'h90;
	   8'h97: op=8'h88;
	   8'h98: op=8'h46;
	   8'h99: op=8'hee;
	   8'h9a: op=8'hb8;
	   8'h9b: op=8'h14;
	   8'h9c: op=8'hde;
	   8'h9d: op=8'h5e;
	   8'h9e: op=8'h0b;
	   8'h9f: op=8'hdb;
	   8'ha0: op=8'he0;
	   8'ha1: op=8'h32;
	   8'ha2: op=8'h3a;
	   8'ha3: op=8'h0a;
	   8'ha4: op=8'h49;
	   8'ha5: op=8'h06;
	   8'ha6: op=8'h24;
	   8'ha7: op=8'h5c;
	   8'ha8: op=8'hc2;
	   8'ha9: op=8'hd3;
	   8'haa: op=8'hac;
	   8'hab: op=8'h62;
	   8'hac: op=8'h91;
	   8'had: op=8'h95;
	   8'hae: op=8'he4;
	   8'haf: op=8'h79;
	   8'hb0: op=8'he7;
	   8'hb1: op=8'hc8;
	   8'hb2: op=8'h37;
	   8'hb3: op=8'h6d;
	   8'hb4: op=8'h8d;
	   8'hb5: op=8'hd5;
	   8'hb6: op=8'h4e;
	   8'hb7: op=8'ha9;
	   8'hb8: op=8'h6c;
	   8'hb9: op=8'h56;
	   8'hba: op=8'hf4;
	   8'hbb: op=8'hea;
	   8'hbc: op=8'h65;
	   8'hbd: op=8'h7a;
	   8'hbe: op=8'hae;
	   8'hbf: op=8'h08;
	   8'hc0: op=8'hba;
	   8'hc1: op=8'h78;
	   8'hc2: op=8'h25;
	   8'hc3: op=8'h2e;
	   8'hc4: op=8'h1c;
	   8'hc5: op=8'ha6;
	   8'hc6: op=8'hb4;
	   8'hc7: op=8'hc6;
	   8'hc8: op=8'he8;
	   8'hc9: op=8'hdd;
	   8'hca: op=8'h74;
	   8'hcb: op=8'h1f;
	   8'hcc: op=8'h4b;
	   8'hcd: op=8'hbd;
	   8'hce: op=8'h8b;
	   8'hcf: op=8'h8a;
	   8'hd0: op=8'h70;
	   8'hd1: op=8'h3e;
	   8'hd2: op=8'hb5;
	   8'hd3: op=8'h66;
	   8'hd4: op=8'h48;
	   8'hd5: op=8'h03;
	   8'hd6: op=8'hf6;
	   8'hd7: op=8'h0e;
	   8'hd8: op=8'h61;
	   8'hd9: op=8'h35;
	   8'hda: op=8'h57;
	   8'hdb: op=8'hb9;
	   8'hdc: op=8'h86;
	   8'hdd: op=8'hc1;
	   8'hde: op=8'h1d;
	   8'hdf: op=8'h9e;
	   8'he0: op=8'he1;
	   8'he1: op=8'hf8;
	   8'he2: op=8'h98;
	   8'he3: op=8'h11;
	   8'he4: op=8'h69;
	   8'he5: op=8'hd9;
	   8'he6: op=8'h8e;
	   8'he7: op=8'h94;
	   8'he8: op=8'h9b;
	   8'he9: op=8'h1e;
	   8'hea: op=8'h87;
	   8'heb: op=8'he9;
	   8'hec: op=8'hce;
	   8'hed: op=8'h55;
	   8'hee: op=8'h28;
	   8'hef: op=8'hdf;
	   8'hf0: op=8'h8c;
	   8'hf1: op=8'ha1;
	   8'hf2: op=8'h89;
	   8'hf3: op=8'h0d;
	   8'hf4: op=8'hbf;
	   8'hf5: op=8'he6;
	   8'hf6: op=8'h42;
	   8'hf7: op=8'h68;
	   8'hf8: op=8'h41;
	   8'hf9: op=8'h99;
	   8'hfa: op=8'h2d;
	   8'hfb: op=8'h0f;
	   8'hfc: op=8'hb0;
	   8'hfd: op=8'h54;
	   8'hfe: op=8'hbb;
	   8'hff: op=8'h16;
	endcase

endmodule




