* /home/sumanto/Desktop/verilog/eSim/transmissiongate/transmissiongate.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Nov  8 20:24:14 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U2-Pad1_ Net-_U2-Pad2_ Net-_U2-Pad3_ jtransmissiongate		
U4  a control Net-_U2-Pad1_ Net-_U2-Pad2_ adc_bridge_2		
v1  a GND pulse		
v2  control GND pulse		
U1  a plot_v1		
U3  control plot_v1		
U6  out plot_v1		
U5  Net-_U2-Pad3_ out dac_bridge_1		

.end
