module m12(output Y, input A, B);
    and(Y, A, B); 
    $dumpvars
endmodule
