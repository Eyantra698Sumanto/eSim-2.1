* /home/sumanto/Desktop/verilog/eSim/boothmultiplier/boothmultiplier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Mon Nov 15 13:14:24 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
v1  Net-_U4-Pad1_ GND pulse		
v2  Net-_U4-Pad2_ GND pulse		
U6  out plot_v1		
U4  Net-_U4-Pad1_ Net-_U4-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U5  Net-_U3-Pad9_ out dac_bridge_1		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ counter4bit		
U2  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ counter4bit		
U3  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U2-Pad3_ Net-_U2-Pad4_ Net-_U2-Pad5_ Net-_U2-Pad6_ Net-_U3-Pad9_ ? ? ? ? ? ? ? jboothmultiplier		

.end
