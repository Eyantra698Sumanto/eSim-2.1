* /home/sumanto/Desktop/verilog/eSim/arraymultiplier/arraymultiplier.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun Nov  7 15:31:20 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U2  Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ Net-_U2-Pad9_ ? ? ? ? ? ? ? junsignedarraymultiplier		
v1  Net-_U5-Pad1_ GND pulse		
v2  Net-_U5-Pad2_ GND pulse		
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ Net-_U1-Pad4_ Net-_U1-Pad5_ Net-_U1-Pad6_ Net-_U1-Pad7_ Net-_U1-Pad8_ Net-_U1-Pad9_ Net-_U1-Pad10_ counter8bit		
U4  out plot_v1		
U5  Net-_U5-Pad1_ Net-_U5-Pad2_ Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
U3  Net-_U2-Pad9_ out dac_bridge_1		

.end
