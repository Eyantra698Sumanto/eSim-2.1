/* verilator lint_off UNUSED */
module jbuffer(a,y);
	input a;
	output y;
	assign y=a;	
endmodule

