* /home/sumanto/Desktop/verilog/eSim/divideby45/divideby45.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Sun Nov 21 16:58:15 2021

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
U1  Net-_U1-Pad1_ Net-_U1-Pad2_ Net-_U1-Pad3_ clk_div_45		
U3  Net-_U1-Pad3_ clkdivideby4_5 dac_bridge_1		
U2  clk en Net-_U1-Pad1_ Net-_U1-Pad2_ adc_bridge_2		
v1  clk GND pulse		
v2  en GND pulse		
U4  clkdivideby4_5 plot_v1		
U5  clk plot_v1		
U6  en plot_v1		

.end
